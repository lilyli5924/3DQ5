library verilog;
use verilog.vl_types.all;
entity experiment2a_v_unit is
end experiment2a_v_unit;
