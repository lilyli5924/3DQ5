library verilog;
use verilog.vl_types.all;
entity tb_experiment4 is
end tb_experiment4;
