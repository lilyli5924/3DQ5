library verilog;
use verilog.vl_types.all;
entity tb_experiment2b_v_unit is
end tb_experiment2b_v_unit;
