library verilog;
use verilog.vl_types.all;
entity tb_experiment1 is
end tb_experiment1;
