library verilog;
use verilog.vl_types.all;
entity experiment2b_v_unit is
end experiment2b_v_unit;
