library verilog;
use verilog.vl_types.all;
entity tb_experiment1_v_unit is
end tb_experiment1_v_unit;
